* SPICE NETLIST
***************************************

.SUBCKT Inverter
** N=4 EP=0 IP=0 FDC=2
M0 3 1 2 nmos L=4.8e-06 W=9.6e-06 AD=1.152e-11 AS=1.152e-11 $X=28800 $Y=-52800 $D=1
M1 4 1 3 pmos L=4.8e-06 W=1.92e-05 AD=2.304e-11 AS=2.304e-11 $X=9600 $Y=24000 $D=0
.ENDS
***************************************
